grammar edu:umn:cs:melt:exts:ableC:libskeleton;

exports edu:umn:cs:melt:exts:ableC:libskeleton:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:libskeleton:concretesyntax;

